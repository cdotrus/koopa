-- Project: {{ koopa.project }}
-- Entity: {{ koopa.name }}


library ieee;
use ieee.std_logic_1164.all;

entity {{ koopa.name }} is 
  generic(

  );
  port(

  );
end entity;


architecture rtl of {{ koopa.name }} is

begin


end architecture;
